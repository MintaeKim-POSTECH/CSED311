`include "macro.v"

module haz_detect_unit (hazard, output_sth, input_sth);
endmodule
